created file






Change on master on github


  This is a change I make on the local master branch, but I want to move it to the remote branch.

    also want to move this to the branch 






Change on branch made on github
















I want this here, and above the things from the branch should be left unharmed
Adding this here on github


do omething on master here
Do one more thing on master here

