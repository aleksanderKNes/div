created file






Change on master on github











Change on branch made on github
