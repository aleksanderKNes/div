created file






Change on master on github


  This is a change I make on the local master branch, but I want to move it to the remote branch.

    also want to move this to the branch 






Change on branch made on github


locally on master

remote on branch made on github



locally on feature

3 Remotely 
4 local, want to move to branch

7, remote commit. AND 8, remote commit


I want this here, and above the things from the branch should be left unharmed
Adding this here on github


do omething on master here
Do one more thing on master here

