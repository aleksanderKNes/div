created file



Writing something on github in a branch created on github
