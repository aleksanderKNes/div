created file






Change on master on github
